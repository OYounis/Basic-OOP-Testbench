package alu_pkg;
`include "random.svh"
`include "coverage.svh"
`include "tester.svh"
`include "scoreboard.svh"
`include "testbench.svh"
endpackage : alu_pkg