class random;
    rand bit [31:0] a;
    rand bit [31:0] b;
    rand bit [2:0] op_code;
endclass
